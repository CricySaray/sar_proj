VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO L28_BOAC_op1_55_6um_stagger_133X74D3
  CLASS COVER ;
  ORIGIN -1.5 -10.5 ;
  FOREIGN L28_BOAC_op1_55_6um_stagger_133X74D3 1.5 10.5 ;
  SIZE 130 BY 62.3 ;
  SYMMETRY X Y ;
  
  OBS
    LAYER ME8 ;
      RECT 0 68.65 133 74.3 ;
      RECT 128 0 133 74.3 ;
      RECT 122 0 125 74.3 ;
      RECT 116 0 119 74.3 ;
      RECT 110 0 113 74.3 ;
      RECT 104 0 107 74.3 ;
      RECT 98 0 101 74.3 ;
      RECT 92 0 95 74.3 ;
      RECT 86 0 89 74.3 ;
      RECT 80 0 83 74.3 ;
      RECT 74 0 77 74.3 ;
      RECT 68 0 71 74.3 ;
      RECT 62 0 65 74.3 ;
      RECT 56 0 59 74.3 ;
      RECT 50 0 53 74.3 ;
      RECT 44 0 47 74.3 ;
      RECT 38 0 41 74.3 ;
      RECT 32 0 35 74.3 ;
      RECT 26 0 29 74.3 ;
      RECT 20 0 23 74.3 ;
      RECT 14 0 17 74.3 ;
      RECT 8 0 11 74.3 ;
      RECT 0 0 5 74.3 ;
      RECT 0 62.65 133 65.65 ;
      RECT 0 56.65 133 59.65 ;
      RECT 0 50.65 133 53.65 ;
      RECT 0 44.65 133 47.65 ;
      RECT 0 38.65 133 41.65 ;
      RECT 0 32.65 133 35.65 ;
      RECT 0 26.65 133 29.65 ;
      RECT 0 20.65 133 23.65 ;
      RECT 0 14.65 133 17.65 ;
      RECT 0 0 133 11.65 ;
    LAYER TMV_RDL ;
      RECT 127.5 0.5 130.5 3.5 ;
      RECT 127.5 5.5 130.5 8.5 ;
      RECT 122.5 0.5 125.5 3.5 ;
      RECT 122.5 5.5 125.5 8.5 ;
      RECT 117.5 0.5 120.5 3.5 ;
      RECT 117.5 5.5 120.5 8.5 ;
      RECT 112.5 0.5 115.5 3.5 ;
      RECT 112.5 5.5 115.5 8.5 ;
      RECT 107.5 0.5 110.5 3.5 ;
      RECT 107.5 5.5 110.5 8.5 ;
      RECT 102.5 0.5 105.5 3.5 ;
      RECT 102.5 5.5 105.5 8.5 ;
      RECT 97.5 0.5 100.5 3.5 ;
      RECT 97.5 5.5 100.5 8.5 ;
      RECT 92.5 0.5 95.5 3.5 ;
      RECT 92.5 5.5 95.5 8.5 ;
      RECT 87.5 0.5 90.5 3.5 ;
      RECT 87.5 5.5 90.5 8.5 ;
      RECT 82.5 0.5 85.5 3.5 ;
      RECT 82.5 5.5 85.5 8.5 ;
      RECT 77.5 0.5 80.5 3.5 ;
      RECT 77.5 5.5 80.5 8.5 ;
      RECT 72.5 0.5 75.5 3.5 ;
      RECT 72.5 5.5 75.5 8.5 ;
      RECT 67.5 0.5 70.5 3.5 ;
      RECT 67.5 5.5 70.5 8.5 ;
      RECT 62.5 0.5 65.5 3.5 ;
      RECT 62.5 5.5 65.5 8.5 ;
      RECT 57.5 0.5 60.5 3.5 ;
      RECT 57.5 5.5 60.5 8.5 ;
      RECT 52.5 0.5 55.5 3.5 ;
      RECT 52.5 5.5 55.5 8.5 ;
      RECT 47.5 0.5 50.5 3.5 ;
      RECT 47.5 5.5 50.5 8.5 ;
      RECT 42.5 0.5 45.5 3.5 ;
      RECT 42.5 5.5 45.5 8.5 ;
      RECT 37.5 0.5 40.5 3.5 ;
      RECT 37.5 5.5 40.5 8.5 ;
      RECT 32.5 0.5 35.5 3.5 ;
      RECT 32.5 5.5 35.5 8.5 ;
      RECT 27.5 0.5 30.5 3.5 ;
      RECT 27.5 5.5 30.5 8.5 ;
      RECT 22.5 0.5 25.5 3.5 ;
      RECT 22.5 5.5 25.5 8.5 ;
      RECT 17.5 0.5 20.5 3.5 ;
      RECT 17.5 5.5 20.5 8.5 ;
      RECT 12.5 0.5 15.5 3.5 ;
      RECT 12.5 5.5 15.5 8.5 ;
      RECT 7.5 0.5 10.5 3.5 ;
      RECT 7.5 5.5 10.5 8.5 ;
      RECT 2.5 0.5 5.5 3.5 ;
      RECT 2.5 5.5 5.5 8.5 ;
    LAYER AL_RDL ;
      RECT 0 0 133 74.3 ;
#    LAYER PASV_RDL ;
#      RECT 1.5 10.5 131.5 72.8 ;
#    LAYER PADMARK ;
#      RECT 0 0 133 74.3 ;
  END
END L28_BOAC_op1_55_6um_stagger_133X74D3

END LIBRARY
