VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO CUT_OSC
  CLASS PAD ;
  ORIGIN 0 0 ;
  FOREIGN CUT_OSC 0 0 ;
  SIZE 90 BY 165 ;
  SYMMETRY X Y R90 ;
  SITE iocore_d ;
  PIN IO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME7 ;
        RECT 31.5 15 61.5 19.5 ;
        RECT 31.5 87.2 61.5 91.7 ;
    END
  END IO
  PIN GNDK
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME7 ;
        RECT 12.5 125.2 90 129.7 ;
        RECT 3.35 141.7 90 146.2 ;
    END
  END GNDK
  PIN GNDI
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME7 ;
        RECT 0 103.6 85.5 106.6 ;
        RECT 4 119.7 85.5 124.2 ;
    END
  END GNDI
  PIN GNDIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME7 ;
        RECT 3.45 3 90.5 7.5 ;
        RECT 3.45 8.5 90.5 13 ;
        RECT 3.45 38.6 90.5 42.5 ;
        RECT 3.45 43.5 90.5 48 ;
        RECT 3.45 49 90.5 51.5 ;
    END
  END GNDIO
  PIN GNDO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME7 ;
        RECT 0 22 87.04 26.5 ;
        RECT 0 27.5 87.04 32 ;
        RECT 0 33 87.04 37.5 ;
        RECT 0 93.1 85.5 95.1 ;
    END
  END GNDO
  OBS
    LAYER ME1 SPACING 0.05 ;
      RECT 0 0 90 165 ;
    LAYER ME2 SPACING 0.05 ;
      RECT 0 0 90 165 ;
    LAYER ME3 SPACING 0.05 ;
      RECT 0 0 90 165 ;
    LAYER ME4 SPACING 0.05 ;
      RECT 0 0 90 165 ;
    LAYER ME5 ;
      RECT 0 93.1 85.51 95.1 ;
      RECT -0.075 93.1 85.51 95.09 ;
      RECT 65.86 3 90.5 7.5 ;
      RECT 65.86 8.5 90.5 13 ;
      RECT 65.86 38.625 90.5 42.5 ;
      RECT 65.86 43.5 90.5 48 ;
      RECT 65.86 49 90.5 51.5 ;
      RECT 65 125.2 90 129.7 ;
      RECT 65 141.7 90 146.2 ;
      RECT 0 103.6 24.06 106.655 ;
      RECT 0 22 20.9 26.5 ;
      RECT 0 27.5 20.9 32 ;
      RECT 0 33 20.9 37.5 ;
      RECT 0 147.6 17 150.6 ;
      RECT 0 151.6 17 154.6 ;
      RECT 0 123.6 8.5 126.6 ;
      RECT 0 127.6 8.5 130.6 ;
      RECT 0 131.6 8.5 134.6 ;
    LAYER ME5 SPACING 0.05 ;
      RECT 0 0 90 165 ;
    LAYER ME6 ;
      RECT 0 93.1 85.5 95.1 ;
      RECT -0.075 93.1 85.505 95.09 ;
      RECT 65.86 3 90.5 7.5 ;
      RECT 65.86 8.5 90.5 13 ;
      RECT 65.86 38.625 90.5 42.5 ;
      RECT 65.86 43.5 90.5 48 ;
      RECT 65.86 49 90.5 51.5 ;
      RECT 65 125.2 90 129.7 ;
      RECT 65 141.7 90 146.2 ;
      RECT 0 103.6 44.96 106.6 ;
      RECT 0 22 20.9 26.5 ;
      RECT 0 27.5 20.9 32 ;
      RECT 0 33 20.9 37.5 ;
      RECT 0 147.6 17 150.6 ;
      RECT 0 151.6 17 154.6 ;
      RECT 0 123.6 8.5 126.6 ;
      RECT 0 127.6 8.5 130.6 ;
      RECT 0 131.6 8.5 134.6 ;
    LAYER ME6 SPACING 0.05 ;
      RECT 0 0 90 165 ;
    LAYER ME7 ;
      RECT 3.45 53.25 85.35 57.75 ;
      RECT 76.38 53 80.78 57.75 ;
      RECT 50.98 53 55.38 57.75 ;
      RECT 30.08 53 34.48 57.75 ;
      RECT 9.15 53 13.55 57.75 ;
      RECT 78.5 147.7 83 154.6 ;
      RECT 67.5 147.7 72 154.6 ;
      RECT 56.5 147.7 61 154.6 ;
      RECT 45.5 147.7 50 154.6 ;
      RECT 34.5 147.7 39 154.6 ;
      RECT 23.5 147.7 28 154.6 ;
      RECT 0 151.6 17 154.6 ;
      RECT 12.5 147.7 17 154.6 ;
      RECT 3.35 147.7 7.85 154.6 ;
      RECT 0 147.7 83 150.6 ;
      RECT 0 147.6 1.85 150.6 ;
      RECT 0 127.6 8.5 130.6 ;
      RECT 4 125.7 8.5 130.6 ;
      RECT 0 125.7 8.5 126.6 ;
      RECT 0 123.6 2.5 126.6 ;
      RECT 81 96.6 85.5 102.1 ;
      RECT 81 108.1 85.5 118.2 ;
      RECT 78.5 131.2 83 140.2 ;
      RECT 75.5 96.6 80 102.1 ;
      RECT 75.5 108.1 80 118.2 ;
      RECT 70 96.6 74.5 102.1 ;
      RECT 70 108.1 74.5 118.2 ;
      RECT 67.5 131.2 72 140.2 ;
      RECT 64.5 96.6 69 102.1 ;
      RECT 64.5 108.1 69 118.2 ;
      RECT 63 87.2 63.5 91.6 ;
      RECT 59 96.6 63.5 102.1 ;
      RECT 59 108.1 63.5 118.2 ;
      RECT 56.5 131.2 61 140.2 ;
      RECT 53.5 96.6 58 102.1 ;
      RECT 53.5 108.1 58 118.2 ;
      RECT 48 96.6 52.5 102.1 ;
      RECT 48 108.1 52.5 118.2 ;
      RECT 45.5 131.2 50 140.2 ;
      RECT 42.5 96.6 47 102.1 ;
      RECT 42.5 108.1 47 118.2 ;
      RECT 37 96.6 41.5 102.1 ;
      RECT 37 108.1 41.5 118.2 ;
      RECT 34.5 131.2 39 140.2 ;
      RECT 31.5 96.6 36 102.1 ;
      RECT 31.5 108.1 36 118.2 ;
      RECT 26 96.6 30.5 102.1 ;
      RECT 26 108.1 30.5 118.2 ;
      RECT 23.5 131.2 28 140.2 ;
      RECT 20.5 96.6 25 102.1 ;
      RECT 20.5 108.1 25 118.2 ;
      RECT 15 96.6 19.5 102.1 ;
      RECT 15 108.1 19.5 118.2 ;
      RECT 12.5 131.2 17 140.2 ;
      RECT 9.5 96.6 14 102.1 ;
      RECT 9.5 108.1 14 118.2 ;
      RECT 4 96.6 8.5 102.1 ;
      RECT 4 108.1 8.5 118.2 ;
      RECT 0 131.6 8.5 134.6 ;
    LAYER ME7 SPACING 0.4 ;
      RECT 87.7 13.66 90 37.94 ;
      RECT 0 20.16 90 21.34 ;
      RECT 62.16 13.66 90 21.34 ;
      RECT 0 13.66 30.84 21.34 ;
      RECT 0 13.66 90 14.34 ;
      RECT 0 0 2.79 21.34 ;
      RECT 0 0 90 2.34 ;
      RECT 0 146.86 90 165 ;
      RECT 0 107.26 2.69 165 ;
      RECT 0 130.36 90 141.04 ;
      RECT 0 124.86 11.84 141.04 ;
      RECT 0 107.26 3.34 141.04 ;
      RECT 86.16 52.16 90 124.54 ;
      RECT 0 107.26 90 119.04 ;
      RECT 0 95.76 90 102.94 ;
      RECT 62.16 52.16 90 92.44 ;
      RECT 0 52.16 30.84 92.44 ;
      RECT 0 52.16 90 86.54 ;
      RECT 0 38.16 2.79 92.44 ;
    LAYER ME8 SPACING 0.4 ;
      RECT 87.7 13.66 90 37.94 ;
      RECT 0 20.16 90 21.34 ;
      RECT 62.16 13.66 90 21.34 ;
      RECT 0 13.66 30.84 21.34 ;
      RECT 0 13.66 90 14.34 ;
      RECT 0 0 2.79 21.34 ;
      RECT 0 0 90 2.34 ;
      RECT 0 146.86 90 165 ;
      RECT 0 107.26 2.69 165 ;
      RECT 0 130.36 90 141.04 ;
      RECT 0 124.86 11.84 141.04 ;
      RECT 0 107.26 3.34 141.04 ;
      RECT 86.16 52.16 90 124.54 ;
      RECT 0 107.26 90 119.04 ;
      RECT 0 95.76 90 102.94 ;
      RECT 62.16 52.16 90 92.44 ;
      RECT 0 52.16 30.84 92.44 ;
      RECT 0 52.16 90 86.54 ;
      RECT 0 38.16 2.79 92.44 ;
  END
END CUT_OSC

END LIBRARY
