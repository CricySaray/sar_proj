VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO L28_BOAC_op1_55_6um_stagger_65D3X74D3
  CLASS COVER ;
  ORIGIN -1.5 -10.5 ;
  FOREIGN L28_BOAC_op1_55_6um_stagger_65D3X74D3 1.5 10.5 ;
  SIZE 62.3 BY 62.3 ;
  SYMMETRY X Y ;

  OBS
    LAYER ME8 ;
      RECT 0 68.65 65.3 74.3 ;
      RECT 61.15 0 65.3 74.3 ;
      RECT 55.15 0 58.15 74.3 ;
      RECT 49.15 0 52.15 74.3 ;
      RECT 43.15 0 46.15 74.3 ;
      RECT 37.15 0 40.15 74.3 ;
      RECT 31.15 0 34.15 74.3 ;
      RECT 25.15 0 28.15 74.3 ;
      RECT 19.15 0 22.15 74.3 ;
      RECT 13.15 0 16.15 74.3 ;
      RECT 7.15 0 10.15 74.3 ;
      RECT 0 0 4.15 74.3 ;
      RECT 0 62.65 65.3 65.65 ;
      RECT 0 56.65 65.3 59.65 ;
      RECT 0 50.65 65.3 53.65 ;
      RECT 0 44.65 65.3 47.65 ;
      RECT 0 38.65 65.3 41.65 ;
      RECT 0 32.65 65.3 35.65 ;
      RECT 0 26.65 65.3 29.65 ;
      RECT 0 20.65 65.3 23.65 ;
      RECT 0 14.65 65.3 17.65 ;
      RECT 0 0 65.3 11.65 ;
    LAYER TMV_RDL ;
      RECT 61.15 0.5 64.15 3.5 ;
      RECT 61.15 5.5 64.15 8.5 ;
      RECT 56.15 0.5 59.15 3.5 ;
      RECT 56.15 5.5 59.15 8.5 ;
      RECT 51.15 0.5 54.15 3.5 ;
      RECT 51.15 5.5 54.15 8.5 ;
      RECT 46.15 0.5 49.15 3.5 ;
      RECT 46.15 5.5 49.15 8.5 ;
      RECT 41.15 0.5 44.15 3.5 ;
      RECT 41.15 5.5 44.15 8.5 ;
      RECT 36.15 0.5 39.15 3.5 ;
      RECT 36.15 5.5 39.15 8.5 ;
      RECT 31.15 0.5 34.15 3.5 ;
      RECT 31.15 5.5 34.15 8.5 ;
      RECT 26.15 0.5 29.15 3.5 ;
      RECT 26.15 5.5 29.15 8.5 ;
      RECT 21.15 0.5 24.15 3.5 ;
      RECT 21.15 5.5 24.15 8.5 ;
      RECT 16.15 0.5 19.15 3.5 ;
      RECT 16.15 5.5 19.15 8.5 ;
      RECT 11.15 0.5 14.15 3.5 ;
      RECT 11.15 5.5 14.15 8.5 ;
      RECT 6.15 0.5 9.15 3.5 ;
      RECT 6.15 5.5 9.15 8.5 ;
      RECT 1.15 0.5 4.15 3.5 ;
      RECT 1.15 5.5 4.15 8.5 ;
    LAYER AL_RDL ;
      RECT 0 0 65.3 74.3 ;
#    LAYER PASV_RDL ;
#      RECT 1.5 10.5 63.8 72.8 ;
#    LAYER PADMARK ;
#      RECT 0 0 65.3 74.3 ;
  END
END L28_BOAC_op1_55_6um_stagger_65D3X74D3

END LIBRARY
