VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO L28_BOAC_op1_55_6um_stagger_picth78_50D8X74D3
  CLASS COVER ;
  ORIGIN -1.5 -10.5 ;
  FOREIGN L28_BOAC_op1_55_6um_stagger_picth78_50D8X74D3 1.5 10.5 ;
  SIZE 47.8 BY 62.3 ;
  SYMMETRY X Y ;
  
  OBS
    LAYER ME7 ;
      RECT 14.4 8 36.4 12.4 ;
    LAYER ME8 ;
      RECT 0 68.65 50.8 74.3 ;
      RECT 44.9 0 50.8 74.3 ;
      RECT 38.9 0 41.9 74.3 ;
      RECT 32.9 0 35.9 74.3 ;
      RECT 26.9 0 29.9 74.3 ;
      RECT 20.9 0 23.9 74.3 ;
      RECT 14.9 0 17.9 74.3 ;
      RECT 8.9 0 11.9 74.3 ;
      RECT 0 0 5.9 74.3 ;
      RECT 0 62.65 50.8 65.65 ;
      RECT 0 56.65 50.8 59.65 ;
      RECT 0 50.65 50.8 53.65 ;
      RECT 0 44.65 50.8 47.65 ;
      RECT 0 38.65 50.8 41.65 ;
      RECT 0 32.65 50.8 35.65 ;
      RECT 0 26.65 50.8 29.65 ;
      RECT 0 20.65 50.8 23.65 ;
      RECT 0 0 50.8 17.65 ;
    LAYER TMV_RDL ;
      RECT 46.4 0.5 49.4 3.5 ;
      RECT 46.4 5.5 49.4 8.5 ;
      RECT 41.4 0.5 44.4 3.5 ;
      RECT 41.4 5.5 44.4 8.5 ;
      RECT 36.4 0.5 39.4 3.5 ;
      RECT 36.4 5.5 39.4 8.5 ;
      RECT 31.4 0.5 34.4 3.5 ;
      RECT 31.4 5.5 34.4 8.5 ;
      RECT 26.4 0.5 29.4 3.5 ;
      RECT 26.4 5.5 29.4 8.5 ;
      RECT 21.4 0.5 24.4 3.5 ;
      RECT 21.4 5.5 24.4 8.5 ;
      RECT 16.4 0.5 19.4 3.5 ;
      RECT 16.4 5.5 19.4 8.5 ;
      RECT 11.4 0.5 14.4 3.5 ;
      RECT 11.4 5.5 14.4 8.5 ;
      RECT 6.4 0.5 9.4 3.5 ;
      RECT 6.4 5.5 9.4 8.5 ;
      RECT 1.4 0.5 4.4 3.5 ;
      RECT 1.4 5.5 4.4 8.5 ;
    LAYER AL_RDL ;
      RECT 0 0 50.8 74.3 ;
#    LAYER PASV_RDL ;
#      RECT 1.5 10.5 49.3 72.8 ;
#    LAYER PADMARK ;
#      RECT 0 0 50.8 74.3 ;
  END
END L28_BOAC_op1_55_6um_stagger_picth78_50D8X74D3

END LIBRARY
