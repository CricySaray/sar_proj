VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO CUTGD
  CLASS ENDCAP BOTTOMLEFT ;
  ORIGIN 0 0 ;
  FOREIGN CUTGD 0 0 ;
  SIZE 50 BY 165 ;
  SYMMETRY X Y R90 ;
  SITE iocore_d ;
  PIN GNDO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME7 ;
        RECT 0 5.5 50 10 ;
        RECT 0 11 50 15.5 ;
        RECT 0 16.5 50 21 ;
        RECT 0 22 50 26.5 ;
        RECT 0 27.5 50 32 ;
        RECT 0 33 50 37.5 ;
        RECT 0 41.275 50 43.275 ;
        RECT 0 93.1 50 95.1 ;
    END
  END GNDO
  PIN GNDI
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME7 ;
        RECT 0 103.6 50 106.6 ;
        RECT 0 127.6 50 130.6 ;
        RECT 0 131.6 50 134.6 ;
    END
  END GNDI
  PIN GNDK
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ME7 ;
        RECT 0 147.6 50 150.6 ;
        RECT 0 151.6 50 154.6 ;
    END
  END GNDK
  OBS
    LAYER ME1 SPACING 0.05 ;
      RECT 0 0 50 165 ;
    LAYER ME2 SPACING 0.05 ;
      RECT 0 0 50 165 ;
    LAYER ME3 SPACING 0.05 ;
      RECT 0 0 50 165 ;
    LAYER ME4 ;
      RECT 0 93.1 50 95.1 ;
      RECT 0 103.6 50 106.6 ;
      RECT 0 127.6 50 130.6 ;
      RECT 0 131.6 50 134.6 ;
      RECT 0 147.6 50 150.6 ;
      RECT 0 151.6 50 154.6 ;
    LAYER ME4 SPACING 0.05 ;
      RECT 0 0 50 165 ;
    LAYER ME5 ;
      RECT 0 5.5 50 10 ;
      RECT 0 11 50 15.5 ;
      RECT 0 16.5 50 21 ;
      RECT 0 22 50 26.5 ;
      RECT 0 27.5 50 32 ;
      RECT 0 33 50 37.5 ;
      RECT 0 41.275 50 43.275 ;
      RECT 0 93.1 50 95.1 ;
      RECT 0 103.6 50 106.6 ;
      RECT 0 127.6 50 130.6 ;
      RECT 0 131.6 50 134.6 ;
      RECT 0 147.6 50 150.6 ;
      RECT 0 151.6 50 154.6 ;
    LAYER ME5 SPACING 0.05 ;
      RECT 0 0 50 165 ;
    LAYER ME6 ;
      RECT 0 5.5 50 10 ;
      RECT 0 11 50 15.5 ;
      RECT 0 16.5 50 21 ;
      RECT 0 22 50 26.5 ;
      RECT 0 27.5 50 32 ;
      RECT 0 33 50 37.5 ;
      RECT 0 41.275 50 43.275 ;
      RECT 0 93.1 50 95.1 ;
      RECT 0 103.6 50 106.6 ;
      RECT 0 127.6 50 130.6 ;
      RECT 0 131.6 50 134.6 ;
      RECT 0 147.6 50 150.6 ;
      RECT 0 151.6 50 154.6 ;
    LAYER ME6 SPACING 0.05 ;
      RECT 0 0 50 165 ;
    LAYER ME7 SPACING 0.4 ;
      RECT 0 0 50 4.84 ;
      RECT 0 38.16 50 40.615 ;
      RECT 0 43.935 50 92.44 ;
      RECT 0 95.76 50 102.94 ;
      RECT 0 107.26 50 126.94 ;
      RECT 0 135.26 50 146.94 ;
      RECT 0 155.26 50 165 ;
    LAYER ME8 SPACING 0.4 ;
      RECT 0 0 50 4.84 ;
      RECT 0 38.16 50 40.615 ;
      RECT 0 43.935 50 92.44 ;
      RECT 0 95.76 50 102.94 ;
      RECT 0 107.26 50 126.94 ;
      RECT 0 135.26 50 146.94 ;
      RECT 0 155.26 50 165 ;
  END
END CUTGD

END LIBRARY
